module controller
	(
	input clk,
	input n_rst,
	input stop_found,
	input start_found,
	input byte_received,
	input ack_prep,
	input check_ack,
	input ack_done,
	input rw_mode,
	input address_match,
	input sda_in,
	output reg rx_enable,
	output reg tx_enable,
	output reg read_enable,
	output reg [1:0] sda_mode,
	output reg load_data
	);
	
	reg tmp_rx_enable;
	reg tmp_tx_enable;
	reg tmp_read_enable;
	reg [1:0] tmp_sda_mode;
	reg tmp_load_data;

	typedef enum bit [3:0] {CHECKADDRESS, WAITADDRESS, SENDNACK, SENDACK, LOADDATA, SENDDATA, STOPDATA, CHECKACK, RECNACK, RECACK,IDLE } state_type;
	state_type state, nextstate;

	always @ (posedge clk, negedge n_rst) begin
		if (n_rst == 1'b0) begin
			state <= IDLE;
			rx_enable <= 1'b0;
			tx_enable <= 1'b0;
			read_enable <= 1'b0;
			sda_mode <= 2'b0;
			load_data <= 1'b0;
		end else begin
			state <= nextstate;
			rx_enable <= tmp_rx_enable;
			tx_enable <= tmp_tx_enable;
			read_enable <= tmp_read_enable;
			sda_mode <= tmp_sda_mode;
			load_data <= tmp_load_data;
		end
	end
	
  always @ (state, stop_found, start_found, byte_received, ack_prep, check_ack, ack_done, rw_mode, address_match, sda_in ) begin : State_Logic
	   nextstate = state;
	   case(state)
	     IDLE: begin
	       if (start_found == 1'b1) begin
	         nextstate = WAITADDRESS;
	       end else begin
	         nextstate = IDLE;
	       end
	     end
	     
	     WAITADDRESS: begin
	       if (ack_prep == 1'b1) begin
	         nextstate = CHECKADDRESS;
	       end else begin
	         nextstate = WAITADDRESS;
	       end
	     end
	     
	     CHECKADDRESS: begin
	       if (address_match == 1'b1 && rw_mode == 1'b1) begin
	         nextstate = SENDACK;
	       end else if (address_match == 1'b0 && rw_mode == 1'b0) begin
	         nextstate = SENDNACK;
	       end else begin
	         nextstate = SENDNACK;
	         //$assert(" Address = 0 and rw mode = 1");
	       end
	     end
	     
	    SENDACK: begin
	      if (check_ack== 1'b1) begin				//was ack_done
	        nextstate = LOADDATA;
	      end else begin
	        nextstate = SENDACK;
	      end
	    end
	    
	    SENDNACK: begin
        if (check_ack == 1'b1) begin			//was ack_done
          nextstate = IDLE;
        end else begin
          nextstate = SENDNACK;
        end
      end
    

    LOADDATA: begin
  
      nextstate = SENDDATA;
      
    end
  

    SENDDATA: begin
      if (byte_received == 1'b1) begin //or ack_prep
        nextstate = STOPDATA;
      end else begin
        nextstate = SENDDATA;
      end
    end

    STOPDATA: begin
      if (ack_prep == 1'b1) begin
        nextstate = CHECKACK;
      end else begin
        nextstate = STOPDATA;
      end
    end


    CHECKACK: begin
      if (check_ack == 1'b1 && sda_in == 1'b0) begin
        nextstate = RECACK;
      end else if (check_ack == 1'b1 && sda_in == 1'b1) begin
        nextstate = RECNACK;
      end
    end


    RECACK: begin
      nextstate = LOADDATA;
    end
    

    RECNACK: begin
      if (stop_found == 1'b1) begin
        nextstate = CHECKADDRESS;
      end else if (stop_found == 1'b0) begin
        nextstate = IDLE;
      end
    end
      
    default: begin
      nextstate = IDLE;
    end
  
  endcase
	end

  always @ (state) begin : Output_Logic
  case(state)

    IDLE: begin
      tmp_rx_enable = 1'b1;
      tmp_tx_enable = 1'b0;
      tmp_read_enable = 1'b0;
      tmp_sda_mode = 2'b00;
      tmp_load_data = 1'b0;
    end
    

    WAITADDRESS: begin
      tmp_rx_enable = 1'b1;
      tmp_tx_enable = 1'b0;
      tmp_read_enable = 1'b0;
      tmp_sda_mode = 2'b00;
      tmp_load_data = 1'b0;
    end
  

    CHECKADDRESS: begin
      tmp_rx_enable = 1'b0;
      tmp_tx_enable = 1'b0;
      tmp_read_enable = 1'b0;
      tmp_sda_mode = 2'b00;
      tmp_load_data = 1'b0;
    end
 

    SENDACK: begin
      tmp_rx_enable = 1'b0;
      tmp_tx_enable = 1'b0;
      tmp_read_enable = 1'b0;
      tmp_sda_mode = 2'b01;
     	tmp_load_data = 1'b0;
    end
 

    SENDNACK: begin
      tmp_rx_enable = 1'b0;
      tmp_tx_enable = 1'b0;
      tmp_read_enable = 1'b0;
      tmp_sda_mode = 2'b10;
      tmp_load_data = 1'b0;
    end
  

    LOADDATA: begin
      tmp_rx_enable = 1'b0;
      tmp_tx_enable = 1'b0;
      tmp_read_enable = 1'b0;
      tmp_sda_mode = 2'b00;
      tmp_load_data = 1'b1;
      
    end
  

    SENDDATA: begin
      tmp_rx_enable = 1'b0;
      tmp_tx_enable = 1'b1;
      tmp_read_enable = 1'b0;
      tmp_sda_mode = 2'b11;
      tmp_load_data = 1'b0;
    end
   
    STOPDATA: begin
      tmp_rx_enable = 1'b0;
      tmp_tx_enable = 1'b0;
      tmp_read_enable = 1'b0;
      tmp_sda_mode = 2'b00;
      tmp_load_data = 1'b0;
    end
    

    CHECKACK: begin
      tmp_rx_enable = 1'b0;
      tmp_tx_enable = 1'b0;
      tmp_read_enable = 1'b0;
      tmp_sda_mode = 2'b00;
      tmp_load_data = 1'b0;
    end

    RECACK: begin
      tmp_rx_enable = 1'b0;
      tmp_tx_enable = 1'b0;
      tmp_read_enable = 1'b1;
      tmp_sda_mode = 2'b00;
      tmp_load_data = 1'b0;
    end
    

    RECNACK: begin
      tmp_rx_enable = 1'b0;
      tmp_tx_enable = 1'b0;
      tmp_read_enable = 1'b0;
      tmp_sda_mode = 2'b00;
      tmp_load_data = 1'b0;
    end
    
    default: begin
      tmp_rx_enable = 1'b1;
      tmp_tx_enable = 1'b0;
      tmp_read_enable = 1'b0;
      tmp_sda_mode = 2'b00;
      tmp_load_data = 1'b0;
    end

  endcase
	end
	
endmodule