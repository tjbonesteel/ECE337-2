module decode
	(
	input wire clk,
	input wire n_rst,
	input wire scl,
	input wire sda_in,
	input wire starting_byte[7:0],
	output wire rw_mode,
	output wire address_match,
	output wire stop_found,
	output wire start_found
	);

	reg scl_1;
	reg scl_2;
	reg sda_1;
	reg sda_2;


	assign address_match = (starting_byte[7:1] && 7'b1111000)? 1'b1 : 1'b0;
	assign start_found = (scl_1 && !scl_2 && sda_1 && sda_2) ? 1'b1 : 1'b0;
	assign stop_found =  (!scl_1 && scl_2 && sda_1 && sda_2) ? 1'b1 : 1'b0;
	assign rw_mode = starting_byte[0];
		
	always @ (posedge clk, negedge n_rst) begin
		if (n_rst == 1'b0) begin
			scl_1 <= 1'b0;
			scl_2 <= 1'b0;
			sda_1 <= 1'b0;
			sda_2 <= 1'b0;
		end else begin
			scl_1 <= scl;
			scl_2 <= scl_1;
			sda_1 <= sda;
			sda_2 <= sda_1;
		end
	end
endmodule
