module avg_four
(
input wire clk,
input wire n_reset,
input wire [15:0] sample_data,
input wire data_ready,
output wire one_k_samples,
output wire modwait,
output wire [15:0] avg_out,
output wire err
);